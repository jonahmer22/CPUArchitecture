module OVERTURE (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_IOSwitch # (.UUID(64'd4 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_0 (.in(wire_1), .en(wire_19), .out(arch_output_value));
  TC_Splitter8 # (.UUID(64'd4503464116114201732 ^ UUID)) Splitter8_1 (.in(wire_2), .out0(wire_29), .out1(wire_4), .out2(wire_13), .out3(wire_6), .out4(wire_28), .out5(wire_16), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd2087377687832881801 ^ UUID)) Decoder3_2 (.dis(wire_23), .sel0(wire_29), .sel1(wire_4), .sel2(wire_13), .out0(wire_12), .out1(wire_30), .out2(wire_18), .out3(wire_21), .out4(wire_26), .out5(wire_31), .out6(wire_19), .out7());
  TC_Decoder3 # (.UUID(64'd686953548377664345 ^ UUID)) Decoder3_3 (.dis(wire_23), .sel0(wire_6), .sel1(wire_28), .sel2(wire_16), .out0(wire_33), .out1(wire_5), .out2(wire_35), .out3(wire_11), .out4(wire_22), .out5(wire_8), .out6(wire_15), .out7());
  TC_Switch # (.UUID(64'd3 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_4 (.en(wire_15), .in(arch_input_value), .out(wire_1_8));
  TC_Not # (.UUID(64'd3770664011524407327 ^ UUID), .BIT_WIDTH(64'd1)) Not_5 (.in(wire_14), .out(wire_23));
  TC_Switch # (.UUID(64'd1759692279329698022 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_6 (.en(wire_14), .in(wire_21), .out(wire_24_0));
  TC_Switch # (.UUID(64'd4057764147882672798 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_7 (.en(wire_0), .in(wire_0), .out(wire_24_1));
  TC_Switch # (.UUID(64'd4197220359267028551 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_8 (.en(wire_0), .in(wire_3), .out(wire_1_2));
  TC_Counter # (.UUID(64'd2126927871900820729 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd1)) Counter8_9 (.clk(clk), .rst(rst), .save(wire_32), .in(wire_17), .out(wire_27));
  TC_Switch # (.UUID(64'd41558568358163725 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_10 (.en(wire_9), .in(wire_9), .out(wire_7_1));
  TC_Switch # (.UUID(64'd4238603235705778763 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_11 (.en(wire_14), .in(wire_12), .out(wire_7_0));
  TC_Switch # (.UUID(64'd2846254507831153103 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_12 (.en(wire_9), .in(wire_2), .out(wire_1_5));
  TC_Switch # (.UUID(64'd3224002108440562466 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_13 (.en(wire_36), .in(wire_25), .out(wire_32));
  TC_Program8_1 # (.UUID(64'd5 ^ UUID), .DEFAULT_FILE_NAME("Program8_1_5.w8.bin"), .ARG_SIG("Program8_1_5=%s")) Program8_1_14 (.clk(clk), .rst(rst), .address(wire_27), .out(wire_2));
  DEC # (.UUID(64'd1943300725040351741 ^ UUID)) DEC_15 (.clk(clk), .rst(rst), .OPCODE(wire_2), .IMMEDIATE(wire_9), .CALCULATION(wire_0), .COPY(wire_14), .CONDITION(wire_36));
  ALU # (.UUID(64'd1628385176953263360 ^ UUID)) ALU_16 (.clk(clk), .rst(rst), .Instruction(wire_2), .Input_1(wire_10), .Input_2(wire_34), .Output(wire_3));
  COND # (.UUID(64'd1052300761800597618 ^ UUID)) COND_17 (.clk(clk), .rst(rst), .Condition(wire_2), .Input(wire_20), .Result(wire_25));
  RegisterPlus # (.UUID(64'd100000 ^ UUID)) RegisterPlus_18 (.clk(clk), .rst(rst), .Load(wire_33), .Save_value(wire_1), .Save(wire_7), .Always_output(wire_17), .Output(wire_1_7));
  RegisterPlus # (.UUID(64'd110000 ^ UUID)) RegisterPlus_19 (.clk(clk), .rst(rst), .Load(wire_5), .Save_value(wire_1), .Save(wire_30), .Always_output(wire_10), .Output(wire_1_4));
  RegisterPlus # (.UUID(64'd120000 ^ UUID)) RegisterPlus_20 (.clk(clk), .rst(rst), .Load(wire_35), .Save_value(wire_1), .Save(wire_18), .Always_output(wire_34), .Output(wire_1_0));
  RegisterPlus # (.UUID(64'd130000 ^ UUID)) RegisterPlus_21 (.clk(clk), .rst(rst), .Load(wire_11), .Save_value(wire_1), .Save(wire_24), .Always_output(wire_20), .Output(wire_1_1));
  RegisterPlus # (.UUID(64'd140000 ^ UUID)) RegisterPlus_22 (.clk(clk), .rst(rst), .Load(wire_22), .Save_value(wire_1), .Save(wire_26), .Always_output(), .Output(wire_1_3));
  RegisterPlus # (.UUID(64'd150000 ^ UUID)) RegisterPlus_23 (.clk(clk), .rst(rst), .Load(wire_8), .Save_value(wire_1), .Save(wire_31), .Always_output(), .Output(wire_1_6));

  wire [0:0] wire_0;
  wire [7:0] wire_1;
  wire [7:0] wire_1_0;
  wire [7:0] wire_1_1;
  wire [7:0] wire_1_2;
  wire [7:0] wire_1_3;
  wire [7:0] wire_1_4;
  wire [7:0] wire_1_5;
  wire [7:0] wire_1_6;
  wire [7:0] wire_1_7;
  wire [7:0] wire_1_8;
  assign wire_1 = wire_1_0|wire_1_1|wire_1_2|wire_1_3|wire_1_4|wire_1_5|wire_1_6|wire_1_7|wire_1_8;
  wire [7:0] wire_2;
  wire [7:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_7_0;
  wire [0:0] wire_7_1;
  assign wire_7 = wire_7_0|wire_7_1;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [7:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  assign arch_input_enable = wire_15;
  wire [0:0] wire_16;
  wire [7:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  assign arch_output_enable = wire_19;
  wire [7:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_24_0;
  wire [0:0] wire_24_1;
  assign wire_24 = wire_24_0|wire_24_1;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [7:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [7:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;

endmodule
