module COND (clk, rst, Condition, Input, Result);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] Condition;
  input  wire [7:0] Input;
  output  wire [0:0] Result;

  TC_Splitter8 # (.UUID(64'd4048989394386344072 ^ UUID)) Splitter8_0 (.in(wire_5), .out0(wire_6), .out1(wire_17), .out2(wire_1), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd1545186655894716180 ^ UUID)) Decoder3_1 (.dis(1'd0), .sel0(wire_6), .sel1(wire_17), .sel2(wire_1), .out0(wire_34), .out1(wire_33), .out2(wire_31), .out3(wire_28), .out4(wire_20), .out5(wire_9), .out6(wire_13), .out7(wire_4));
  TC_Splitter8 # (.UUID(64'd3247615531470452602 ^ UUID)) Splitter8_2 (.in(wire_22), .out0(wire_29), .out1(wire_37), .out2(wire_11), .out3(wire_35), .out4(wire_24), .out5(wire_15), .out6(wire_7), .out7(wire_2));
  TC_And # (.UUID(64'd3266331449444073027 ^ UUID), .BIT_WIDTH(64'd1)) And_3 (.in0(wire_31), .in1(wire_2), .out(wire_21));
  TC_Not # (.UUID(64'd1682344307092799045 ^ UUID), .BIT_WIDTH(64'd1)) Not_4 (.in(wire_34), .out(wire_23));
  TC_Switch # (.UUID(64'd4064409333541083717 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_5 (.en(wire_23), .in(wire_10), .out(wire_14));
  TC_Or3 # (.UUID(64'd717636221321199949 ^ UUID), .BIT_WIDTH(64'd1)) Or3_6 (.in0(wire_29), .in1(wire_37), .in2(wire_11), .out(wire_32));
  TC_Or3 # (.UUID(64'd2919027784872788916 ^ UUID), .BIT_WIDTH(64'd1)) Or3_7 (.in0(wire_32), .in1(wire_35), .in2(wire_24), .out(wire_19));
  TC_Or3 # (.UUID(64'd1055443418004554436 ^ UUID), .BIT_WIDTH(64'd1)) Or3_8 (.in0(wire_19), .in1(wire_15), .in2(wire_7), .out(wire_36));
  TC_Or # (.UUID(64'd3960558216836422499 ^ UUID), .BIT_WIDTH(64'd1)) Or_9 (.in0(wire_36), .in1(wire_2), .out(wire_3));
  TC_Not # (.UUID(64'd3215456452341280849 ^ UUID), .BIT_WIDTH(64'd1)) Not_10 (.in(wire_3), .out(wire_25));
  TC_And # (.UUID(64'd2101890364078172225 ^ UUID), .BIT_WIDTH(64'd1)) And_11 (.in0(wire_33), .in1(wire_25), .out(wire_12));
  TC_Switch # (.UUID(64'd3248473676661519162 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_12 (.en(wire_20), .in(wire_20), .out(wire_10_6));
  TC_Switch # (.UUID(64'd806757236731844138 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_13 (.en(wire_21), .in(wire_21), .out(wire_10_3));
  TC_Switch # (.UUID(64'd75066545321735865 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_14 (.en(wire_12), .in(wire_12), .out(wire_10_0));
  TC_Or # (.UUID(64'd3102264118142632147 ^ UUID), .BIT_WIDTH(64'd1)) Or_15 (.in0(wire_25), .in1(wire_2), .out(wire_26));
  TC_And # (.UUID(64'd3058654970275571168 ^ UUID), .BIT_WIDTH(64'd1)) And_16 (.in0(wire_28), .in1(wire_26), .out(wire_0));
  TC_Switch # (.UUID(64'd3355416313250400733 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_17 (.en(wire_0), .in(wire_0), .out(wire_10_5));
  TC_And # (.UUID(64'd265441578866667544 ^ UUID), .BIT_WIDTH(64'd1)) And_18 (.in0(wire_9), .in1(wire_3), .out(wire_27));
  TC_Switch # (.UUID(64'd1211468010913970906 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_19 (.en(wire_27), .in(wire_27), .out(wire_10_4));
  TC_Not # (.UUID(64'd2332248486572952950 ^ UUID), .BIT_WIDTH(64'd1)) Not_20 (.in(wire_2), .out(wire_30));
  TC_Switch # (.UUID(64'd2721636531639673806 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_21 (.en(wire_16), .in(wire_16), .out(wire_10_1));
  TC_And # (.UUID(64'd2709005807656095038 ^ UUID), .BIT_WIDTH(64'd1)) And_22 (.in0(wire_13), .in1(wire_30), .out(wire_16));
  TC_And3 # (.UUID(64'd2516764302339524543 ^ UUID), .BIT_WIDTH(64'd1)) And3_23 (.in0(wire_4), .in1(wire_3), .in2(wire_18), .out(wire_8));
  TC_Not # (.UUID(64'd2398651143589734285 ^ UUID), .BIT_WIDTH(64'd1)) Not_24 (.in(wire_2), .out(wire_18));
  TC_Switch # (.UUID(64'd3282149085299710672 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_25 (.en(wire_8), .in(wire_8), .out(wire_10_2));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [7:0] wire_5;
  assign wire_5 = Condition;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_10_0;
  wire [0:0] wire_10_1;
  wire [0:0] wire_10_2;
  wire [0:0] wire_10_3;
  wire [0:0] wire_10_4;
  wire [0:0] wire_10_5;
  wire [0:0] wire_10_6;
  assign wire_10 = wire_10_0|wire_10_1|wire_10_2|wire_10_3|wire_10_4|wire_10_5|wire_10_6;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  assign Result = wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [7:0] wire_22;
  assign wire_22 = Input;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;

endmodule
